module And(InA, InB, Out);
    input InA, InB;
    output Out;
    
    assign Out = InA & InB;
endmodule